`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
//
// HUST Verilog Experiment 2.3 - decoder 3 to 8
//
// Pan Yue
//
//////////////////////////////////////////////////////////////////////////////////


module decoder_3to8(in, out);
    input [2:0] in;
    output reg [7:0] out;
    
    always@(in)  
        case(in)  
            3'b000 : out[7:0] = 8'b11111110;
            3'b001 : out[7:0] = 8'b11111101;
            3'b010 : out[7:0] = 8'b11111011;
            3'b011 : out[7:0] = 8'b11110111;
            3'b100 : out[7:0] = 8'b11101111;
            3'b101 : out[7:0] = 8'b11011111;
            3'b110 : out[7:0] = 8'b10111111;
            default : out[7:0] = 8'b01111111;
        endcase
endmodule